interface uart_if;
	logic tx;
	logic rx;
	logic baud_o;
endinterface
